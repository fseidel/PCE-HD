`default_nettype none

/*
 * HuC6270 Verilog Module for Priority Circuit
 *
 * (C) 2018 Ford Seidel and Amolak Nagi
 */

module PriorityCircuit();

endmodule: PriorityCircuit
