`default_nettype none

/*
 * HuC6270 Verilog Module for Receiving sync signals
 *
 * (C) 2018 Ford Seidel and Amolak Nagi
 */

module Sync(input logic clock,
                        HSYNC_n,
                        VSYNC_n);

endmodule: Sync
