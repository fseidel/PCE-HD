`default_nettype none

/*
 * verilog model of HuC6270 VDC Address Unit
 *
 * (C) 2018 Ford Seidel and Amolak Nagi
 */

module AddressUnit (input clock,
                    output logic [15:0] MA // Address signals to VRAM
                    );



endmodule: AddressUnit
